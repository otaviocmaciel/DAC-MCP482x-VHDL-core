LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL; 

entity mcpdactest is
PORT(
    clk     : IN     STD_LOGIC;                             --system clock
    cs	    : OUT    STD_logic;										--chip select
    sclk    : OUT    STD_LOGIC;                             --spi clock
    mosi    : OUT    STD_LOGIC;                             --master out slave in
	SW : IN STD_LOGIC
);
end mcpdactest;

architecture hardware of mcpdactest is

COMPONENT spi
    	PORT(
        	clk 		: IN  STD_LOGIC;
        	reset_n 	: IN  STD_LOGIC;
        	enable 		: IN  STD_LOGIC;
			cpol    	: IN  STD_LOGIC;
			cpha    	: IN  STD_LOGIC;
			miso		: IN  STD_LOGIC;
        	sclk 		: OUT STD_LOGIC;
        	ss_n 		: OUT STD_LOGIC;
        	mosi 		: OUT STD_LOGIC;
        	busy 		: OUT STD_LOGIC;
        	tx 		: IN  STD_LOGIC_VECTOR(15 downto 0);
        	rx 		: OUT STD_LOGIC_VECTOR(15 downto 0)
       		);
END COMPONENT;

-- SPI Signals
SIGNAL TX : STD_LOGIC_VECTOR(15 downto 0);
SIGNAL ENABLE : std_logic;
SIGNAL RX_ENABLE : std_logic := '1';
SIGNAL BUSY : std_logic;
SIGNAL reset_n : std_logic := '0';
SIGNAL rx_master, rx_slave: STD_LOGIC_VECTOR(15 downto 0);
SIGNAL CPHA :STD_LOGIC := '0';
SIGNAL CPOL :STD_LOGIC := '0';
SIGNAL MISO : std_logic;

-- Controls MCP DAC Signals
SIGNAL txA		: STD_LOGIC_VECTOR(11 DOWNTO 0) := "100010111010";
SIGNAL txB		: STD_LOGIC_VECTOR(11 DOWNTO 0) := "101010101010";
SIGNAL DACSel	: STD_LOGIC	:= '0';
SIGNAL DACGain	: STD_LOGIC := '1';
SIGNAL SHDN		: STD_LOGIC := '1';
SIGNAL START 	: STD_LOGIC;

SIGNAL BufferTX 		: STD_LOGIC_VECTOR(15 downto 0);
SIGNAL LastTX_A 	 	: STD_LOGIC_VECTOR(11 downto 0);
SIGNAL LastTX_B 	 	: STD_LOGIC_VECTOR(11 downto 0);
TYPE StateMachine_DAC is (IDLE, TRANSMIT, WAITING);
SIGNAL State_DAC 		: StateMachine_DAC;

-- Sin function array
    type sine_wave_array is array (0 to 359) of std_logic_vector(11 downto 0);
    constant sine_wave : sine_wave_array := (
	 "100000000000", "100000100100", "100001001000", "100001101011", "100010001111", "100010110011", 
	 "100011010111", "100011111010", "100100011110", "100101000001", "100101100100", "100110001000", 
	 "100110101011", "100111001110", "100111110001", "101000010011", "101000110110", "101001011000", 
	 "101001111010", "101010011100", "101010111110", "101011100000", "101100000001", "101100100010", 
	 "101101000011", "101101100011", "101110000100", "101110100100", "101111000011", "101111100011", 
	 "110000000010", "110000100001", "110000111111", "110001011110", "110001111011", "110010011001", 
	 "110010110110", "110011010011", "110011101111", "110100001011", "110100100111", "110101000010", 
	 "110101011101", "110101110111", "110110010001", "110110101011", "110111000100", "110111011100", 
	 "110111110100", "111000001100", "111000100011", "111000111010", "111001010000", "111001100110", 
	 "111001111011", "111010010000", "111010100100", "111010111000", "111011001011", "111011011110", 
	 "111011110000", "111100000001", "111100010010", "111100100011", "111100110011", "111101000010", 
	 "111101010001", "111101011111", "111101101100", "111101111001", "111110000110", "111110010010", 
	 "111110011101", "111110101000", "111110110010", "111110111011", "111111000100", "111111001100", 
	 "111111010100", "111111011011", "111111100001", "111111100111", "111111101100", "111111110001", 
	 "111111110101", "111111111000", "111111111011", "111111111101", "111111111110", "111111111111", 
	 "111111111111", "111111111111", "111111111101", "111111111100", "111111111001", "111111110110", 
	 "111111110011", "111111101111", "111111101010", "111111100100", "111111011110", "111111010111", 
	 "111111010000", "111111001000", "111111000000", "111110110111", "111110101101", "111110100010", 
	 "111110010111", "111110001100", "111110000000", "111101110011", "111101100110", "111101011000", 
	 "111101001001", "111100111010", "111100101011", "111100011011", "111100001010", "111011111001", 
	 "111011100111", "111011010100", "111011000001", "111010101110", "111010011010", "111010000110", 
	 "111001110001", "111001011011", "111001000101", "111000101111", "111000011000", "111000000000", 
	 "110111101000", "110111010000", "110110110111", "110110011110", "110110000100", "110101101010", 
	 "110101001111", "110100110100", "110100011001", "110011111101", "110011100001", "110011000101", 
	 "110010101000", "110010001010", "110001101101", "110001001111", "110000110000", "110000010010", 
	 "101111110011", "101111010011", "101110110100", "101110010100", "101101110100", "101101010011", 
	 "101100110010", "101100010001", "101011110000", "101011001111", "101010101101", "101010001011", 
	 "101001101001", "101001000111", "101000100101", "101000000010", "100111011111", "100110111100", 
	 "100110011001", "100101110110", "100101010011", "100100101111", "100100001100", "100011101000", 
	 "100011000101", "100010100001", "100001111101", "100001011010", "100000110110", "100000010010", 
	 "011111101110", "011111001010", "011110100110", "011110000011", "011101011111", "011100111011", 
	 "011100011000", "011011110100", "011011010001", "011010101101", "011010001010", "011001100111", 
	 "011001000100", "011000100001", "010111111110", "010111011011", "010110111001", "010110010111", 
	 "010101110101", "010101010011", "010100110001", "010100010000", "010011101111", "010011001110", 
	 "010010101101", "010010001100", "010001101100", "010001001100", "010000101101", "010000001101", 
	 "001111101110", "001111010000", "001110110001", "001110010011", "001101110110", "001101011000",
	 "001100111011", "001100011111", "001100000011", "001011100111", "001011001100", "001010110001",
	 "001010010110", "001001111100", "001001100010", "001001001001", "001000110000", "001000011000",
	 "001000000000", "000111101000", "000111010001", "000110111011", "000110100101", "000110001111",
	 "000101111010", "000101100110", "000101010010", "000100111111", "000100101100", "000100011001",
	 "000100000111", "000011110110", "000011100101", "000011010101", "000011000110", "000010110111",
	 "000010101000", "000010011010", "000010001101", "000010000000", "000001110100", "000001101001",
	 "000001011110", "000001010011", "000001001001", "000001000000", "000000111000", "000000110000",
	 "000000101001", "000000100010", "000000011100", "000000010110", "000000010001", "000000001101",
	 "000000001010", "000000000111", "000000000100", "000000000011", "000000000001", "000000000001",
	 "000000000001", "000000000010", "000000000011", "000000000101", "000000001000", "000000001011",
	 "000000001111", "000000010100", "000000011001", "000000011111", "000000100101", "000000101100",
	 "000000110100", "000000111100", "000001000101", "000001001110", "000001011000", "000001100011",
	 "000001101110", "000001111010", "000010000111", "000010010100", "000010100001", "000010101111",
	 "000010111110", "000011001101", "000011011101", "000011101110", "000011111111", "000100010000",
	 "000100100010", "000100110101", "000101001000", "000101011100", "000101110000", "000110000101",
	 "000110011010", "000110110000", "000111000110", "000111011101", "000111110100", "001000001100",
	 "001000100100", "001000111100", "001001010101", "001001101111", "001010001001", "001010100011",
	 "001010111110", "001011011001", "001011110101", "001100010001", "001100101101", "001101001010",
	 "001101100111", "001110000101", "001110100010", "001111000001", "001111011111", "001111111110",
	 "010000011101", "010000111101", "010001011100", "010001111100", "010010011101", "010010111101",
	 "010011011110", "010011111111", "010100100000", "010101000010", "010101100100", "010110000110",
	 "010110101000", "010111001010", "010111101101", "011000001111", "011000110010", "011001010101",
	 "011001111000", "011010011100", "011010111111", "011011100010", "011100000110", "011100101001",
	 "011101001101", "011101110001", "011110010101", "011110111000", "011111011100", "100000000000" 
	 );

    signal index_sin 	: integer range 0 to 359 := 0;
	 signal index_cos 	: integer range 0 to 359 := 90;
	 signal clk_counter 	: integer range 0 to 138 := 0;
	 signal CLK_2			: std_logic := '0'; -- (50MHz/2) -> 25MHz Signal to use in SPI Core
	 
begin
START <= not SW;

process(CLK)
begin
if(falling_edge(CLK)) then
	if clk_counter = 138 then  				-- 138 -> each 2.78 us update the counter
		clk_counter <= 0;
      index_sin <= (index_sin + 1) mod 360; -- 1 steps 
		index_cos <= (index_cos + 1) mod 360; -- 1 step
   else
      clk_counter <= clk_counter + 1;
   end if;
	CLK_2 <= not CLK_2;
end if;
end process;

process(CLK)
begin
if(falling_edge(CLK)) then
	CASE State_DAC is

		When IDLE =>
			reset_n <= '0';
			txA <= sine_wave(index_sin);
			txB <= sine_wave(index_cos);
		
			if(START = '1') then
				if(DACSel = '0' and LastTX_A /= txA) then
					LastTX_A <= txA;
					BufferTX <= '0' & '0' & DACGain & SHDN & txA;
					DACSel <= '1';
					State_DAC <= TRANSMIT;
				elsif(DACSel = '1' and LastTX_B /= txB) then
					LastTX_B <= txB;
					BufferTX <= '1' & '0' & DACGain & SHDN & txB;
					DACSel <= '0';
					State_DAC <= TRANSMIT;
				end if;
			end if;
		
		When TRANSMIT =>
			reset_n <= '1';
			TX <= BufferTX;
			ENABLE <= '1';
			if(BUSY = '1') then
				State_DAC <= WAITING;
			end if;

		When WAITING =>
			if(BUSY = '0') then
				State_DAC <= IDLE;
			end if;

	END CASE;
end if;
end process;

SPI1 : spi port map(
       		clk		=> CLK_2, -- 25MHz to SPI core
        	reset_n		=> reset_n,
        	enable 		=> ENABLE,
		cpol    	=> CPOL,
		cpha    	=> CPHA,
		miso		=> MISO,
        	sclk 		=> sclk,
        	ss_n 		=> cs,
        	mosi 		=> mosi,
        	busy 		=> BUSY,
        	tx 		=> TX,
        	rx 		=> open
);
end hardware;
